`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 07/24/2025 05:42:10 PM
// Design Name: 
// Module Name: divider64
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module divider64 (
    input logic clk_i,
    input logic reset_i,
    input logic stall_i,
    input logic sign_i,
    input logic start_i,
    input logic [63:0] dividend_i, 
    input logic [63:0] divider_i,
    
    output logic [63:0] quotient_o, 
    output logic [63:0] remainder_o,
    output logic valid_o
);
    
    // Internal registers
    logic [63:0] N, D;
    logic [63:0] Q, R;
    logic [63:0] N_r, D_r;
    
    // Control signals
    logic [6:0] n;  // 7 bits to count up to 64
    logic [6:0] bits;
    logic loaded;
    logic N_bit;
    
    // Status signals
    wire logic ready = !n;
    wire logic neg_out;
    wire logic n_sign = dividend_i[63];
    wire logic d_sign = divider_i[63];
    wire logic [63:0] abs_dividend;
    wire logic divide_by_zero;
    wire logic signed_ovf;

    // Output sign calculation
    assign neg_out = sign_i & ((D_r[63] & ~N_r[63]) | (~D_r[63] & N_r[63]));
    
    // Absolute value calculation
    assign abs_dividend = (~(sign_i & n_sign)) ? dividend_i : ~dividend_i + 1'b1;

    // Error conditions
    assign divide_by_zero = loaded && (D_r == 0);
    assign signed_ovf = loaded && sign_i && (N_r == -64'h8000000000000000) && (D_r == -1);
    
    // Bit-width calculation
    always_comb begin
        N_bit = N[n-1'b1];
        if(divide_by_zero || signed_ovf)
            bits = 7'd3;
        else
            casez (abs_dividend)
                64'b0000000000000000000000000000000000000000000000000000000000000001: bits = 7'd3;
                64'b000000000000000000000000000000000000000000000000000000000000001?: bits = 7'd3;
                64'b00000000000000000000000000000000000000000000000000000000000001??: bits = 7'd3;
                64'b0000000000000000000000000000000000000000000000000000000000001???: bits = 7'd4;
                64'b000000000000000000000000000000000000000000000000000000000001????: bits = 7'd5;
                64'b00000000000000000000000000000000000000000000000000000000001?????: bits = 7'd6;
                64'b0000000000000000000000000000000000000000000000000000000001??????: bits = 7'd7;
                64'b000000000000000000000000000000000000000000000000000000001???????: bits = 7'd8;
                64'b00000000000000000000000000000000000000000000000000000001????????: bits = 7'd9;
                64'b0000000000000000000000000000000000000000000000000000001?????????: bits = 7'd10;
                64'b000000000000000000000000000000000000000000000000000001??????????: bits = 7'd11;
                64'b00000000000000000000000000000000000000000000000000001???????????: bits = 7'd12;
                64'b0000000000000000000000000000000000000000000000000001????????????: bits = 7'd13;
                64'b000000000000000000000000000000000000000000000000001?????????????: bits = 7'd14;
                64'b00000000000000000000000000000000000000000000000001??????????????: bits = 7'd15;
                64'b0000000000000000000000000000000000000000000000001???????????????: bits = 7'd16;
                64'b000000000000000000000000000000000000000000000001????????????????: bits = 7'd17;
                64'b00000000000000000000000000000000000000000000001?????????????????: bits = 7'd18;
                64'b0000000000000000000000000000000000000000000001??????????????????: bits = 7'd19;
                64'b000000000000000000000000000000000000000000001???????????????????: bits = 7'd20;
                64'b00000000000000000000000000000000000000000001????????????????????: bits = 7'd21;
                64'b0000000000000000000000000000000000000000001?????????????????????: bits = 7'd22;
                64'b000000000000000000000000000000000000000001??????????????????????: bits = 7'd23;
                64'b00000000000000000000000000000000000000001???????????????????????: bits = 7'd24;
                64'b0000000000000000000000000000000000000001????????????????????????: bits = 7'd25;
                64'b000000000000000000000000000000000000001?????????????????????????: bits = 7'd26;
                64'b00000000000000000000000000000000000001??????????????????????????: bits = 7'd27;
                64'b0000000000000000000000000000000000001???????????????????????????: bits = 7'd28;
                64'b000000000000000000000000000000000001????????????????????????????: bits = 7'd29;
                64'b00000000000000000000000000000000001?????????????????????????????: bits = 7'd30;
                64'b0000000000000000000000000000000001??????????????????????????????: bits = 7'd31;
                64'b000000000000000000000000000000001???????????????????????????????: bits = 7'd32;
                64'b00000000000000000000000000000001????????????????????????????????: bits = 7'd33;
                64'b0000000000000000000000000000001?????????????????????????????????: bits = 7'd34;
                64'b000000000000000000000000000001??????????????????????????????????: bits = 7'd35;
                64'b00000000000000000000000000001???????????????????????????????????: bits = 7'd36;
                64'b0000000000000000000000000001????????????????????????????????????: bits = 7'd37;
                64'b000000000000000000000000001?????????????????????????????????????: bits = 7'd38;
                64'b00000000000000000000000001??????????????????????????????????????: bits = 7'd39;
                64'b0000000000000000000000001???????????????????????????????????????: bits = 7'd40;
                64'b000000000000000000000001????????????????????????????????????????: bits = 7'd41;
                64'b00000000000000000000001?????????????????????????????????????????: bits = 7'd42;
                64'b0000000000000000000001??????????????????????????????????????????: bits = 7'd43;
                64'b000000000000000000001???????????????????????????????????????????: bits = 7'd44;
                64'b00000000000000000001????????????????????????????????????????????: bits = 7'd45;
                64'b0000000000000000001?????????????????????????????????????????????: bits = 7'd46;
                64'b000000000000000001??????????????????????????????????????????????: bits = 7'd47;
                64'b00000000000000001???????????????????????????????????????????????: bits = 7'd48;
                64'b0000000000000001????????????????????????????????????????????????: bits = 7'd49;
                64'b000000000000001?????????????????????????????????????????????????: bits = 7'd50;
                64'b00000000000001??????????????????????????????????????????????????: bits = 7'd51;
                64'b0000000000001???????????????????????????????????????????????????: bits = 7'd52;
                64'b000000000001????????????????????????????????????????????????????: bits = 7'd53;
                64'b00000000001?????????????????????????????????????????????????????: bits = 7'd54;
                64'b0000000001??????????????????????????????????????????????????????: bits = 7'd55;
                64'b000000001???????????????????????????????????????????????????????: bits = 7'd56;
                64'b00000001????????????????????????????????????????????????????????: bits = 7'd57;
                64'b0000001?????????????????????????????????????????????????????????: bits = 7'd58;
                64'b000001??????????????????????????????????????????????????????????: bits = 7'd59;
                64'b00001???????????????????????????????????????????????????????????: bits = 7'd60;
                64'b0001????????????????????????????????????????????????????????????: bits = 7'd61;
                64'b001?????????????????????????????????????????????????????????????: bits = 7'd62;
                64'b01??????????????????????????????????????????????????????????????: bits = 7'd63;
                64'b1???????????????????????????????????????????????????????????????: bits = 7'd64;
                default: bits = 7'd3;
            endcase
    end
    
    // Division algorithm
    wire logic [63:0] r_shift = {R[62:0], N_bit};
    wire logic [63:0] r_diff = (r_shift >= D) ? r_shift - D : r_shift;
    wire logic [63:0] q = (r_shift >= D) ? (1 << (n-1'b1)) : 0;
    
    // Main FSM
    always_ff @(posedge clk_i or negedge reset_i) begin
        if (!reset_i) begin
            n <= 0;
            Q <= 0;
            R <= 0;
            N <= 0;
            D <= 0;
            N_r <= 0;
            D_r <= 0;
            loaded <= 1'b0;
        end
        else if (~stall_i) begin
            // Case 1: Start new division when start_i is asserted and divider is idle
            if (start_i && ready) begin
                n     <= bits;
                Q     <= 0;
                R     <= 0;
                N     <= (~(sign_i & n_sign)) ? dividend_i : ~dividend_i + 1'b1;
                D     <= (~(sign_i & d_sign)) ? divider_i : ~divider_i + 1'b1;
                N_r   <= dividend_i;
                D_r   <= divider_i;
                loaded <= 1'b1;
            end
            // Case 2: Continue division cycle if not finished
            else if (n > 0 && loaded) begin
                n <= n - 1'b1;
                R <= r_diff;
                Q <= Q | q;
            end
            // Case 3: Reset `loaded` once complete and ready for next start
            else if (ready) begin
                loaded <= 1'b0;
            end
        end
    end

    
    // Output generation
    always_comb begin
        if(divide_by_zero) begin
            quotient_o = sign_i ? -1 : 64'hFFFFFFFFFFFFFFFF;
            remainder_o = N_r;
        end
        else if(signed_ovf) begin
            quotient_o = -64'h8000000000000000;
            remainder_o = 0;
        end
        else begin
            quotient_o = (~neg_out) ? Q : ~Q + 1'b1;
            remainder_o = (~(sign_i & N_r[63])) ? R : ~R + 1'b1;
        end
    end
    
    assign valid_o = ready;

endmodule
